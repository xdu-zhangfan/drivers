module spi_com (
    
);
    
endmodule